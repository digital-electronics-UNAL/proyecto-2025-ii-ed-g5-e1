module code #(
   
)(
    input [3:0] digdec,
    output [3:0] dighex
);
endmodule