module LCD1602_controller #(parameter NUM_COMMANDS = 4, 
                                      NUM_DATA_ALL = 32,  
                                      NUM_DATA_PERLINE = 16,
                                      DATA_BITS = 8,
                                      COUNT_MAX = 800000)(
    input clk,            
    input reset,          
    input ready_i,
    output reg rs,     // si lo que llega a la LCD es dato o comando(si es de derecha a izquierda, cursor parpadenate o no)   
    output reg rw,
    output enable,    
    output reg [DATA_BITS-1:0] data
);

// 16-20 Definir los estados de la FSM, param local: acceder desde afuera
localparam IDLE = 3'b000;
localparam CONFIG_CMD1 = 3'b001;
localparam WR_STATIC_TEXT_1L = 3'b010;
localparam CONFIG_CMD2 = 3'b011;
localparam WR_STATIC_TEXT_2L = 3'b100;

reg [2:0] fsm_state;//el estado presente. el que va a saltar entre los valores de localparam
reg [2:0] next_state;
reg clk_16ms;//asiganr la salida enable 

// Comandos de configuración, no van a ser estados de la maquina. SOlo configuraciones del lcd
localparam CLEAR_DISPLAY = 8'h01;
localparam SHIFT_CURSOR_RIGHT = 8'h06;
localparam DISPON_CURSOROFF = 8'h0C;//o uno
localparam DISPON_CURSORBLINK = 8'h0E;//o  el otro
localparam LINES2_MATRIX5x8_MODE8bit = 8'h38; //LD con varios modos. 8 bits al tiempo:en paralelo, O pseudo paralelo usa 4 bits
localparam START_2LINE = 8'hC0; //para arrancar en la segunda linea

//un caracter necesita los 8 bits por D0 a D7
//poder con solo4 bits, con el otro modo, 


// Definir un contador para el divisor de frecuencia
reg [$clog2(COUNT_MAX)-1:0] clk_counter;
// Definir un contador para controlar el envío de comandos
reg [$clog2(NUM_COMMANDS):0] command_counter;
// Definir un contador para controlar el envío de datos
reg [$clog2(NUM_DATA_PERLINE):0] data_counter;

// Banco de registros, como se contruye una memoria, guarda comandos de config
reg [DATA_BITS-1:0] static_data_mem [0: NUM_DATA_ALL-1];//
reg [DATA_BITS-1:0] config_mem [0:NUM_COMMANDS-1]; 

initial begin
    fsm_state <= IDLE;
    command_counter <= 'b0;
    data_counter <= 'b0;
    rs <= 1'b0;
    rw <= 1'b0;
    data <= 8'b0;
    clk_16ms <= 1'b0;
    clk_counter <= 'b0;
    $readmemh("/home/alejandro/github-classroom/digital-electronics-UNAL/lab07-lcd-en-modo-paralelo-2025-ii-ed-g5-e1/src/data.txt", static_data_mem);    //leer txt y llenar memoria
	config_mem[0] <= LINES2_MATRIX5x8_MODE8bit;
	config_mem[1] <= SHIFT_CURSOR_RIGHT;
	config_mem[2] <= DISPON_CURSOROFF;
	config_mem[3] <= CLEAR_DISPLAY;
end

always @(posedge clk) begin
    if (clk_counter == COUNT_MAX-1) begin
        clk_16ms <= ~clk_16ms;
        clk_counter <= 'b0;
    end else begin
        clk_counter <= clk_counter + 1;
    end
end


always @(posedge clk_16ms)begin
    if(reset == 0)begin //logica negada en la FPGA
        fsm_state <= IDLE;
    end else begin
        fsm_state <= next_state;
    end
end

always @(*) begin
    case(fsm_state)
        IDLE: begin //estado inicial
            next_state <= (ready_i)? CONFIG_CMD1 : IDLE;
        end
        CONFIG_CMD1: begin 
            next_state <= (command_counter == NUM_COMMANDS)? WR_STATIC_TEXT_1L : CONFIG_CMD1;
        end
        WR_STATIC_TEXT_1L:begin
			next_state <= (data_counter == NUM_DATA_PERLINE)? CONFIG_CMD2 : WR_STATIC_TEXT_1L;
        end
        CONFIG_CMD2: begin 
            next_state <= WR_STATIC_TEXT_2L;
        end
		WR_STATIC_TEXT_2L: begin
			next_state <= (data_counter == NUM_DATA_PERLINE)? IDLE : WR_STATIC_TEXT_2L;
		end
        default: next_state = IDLE;
    endcase
end

always @(posedge clk_16ms) begin
    if (reset == 0) begin
        command_counter <= 'b0;
        data_counter <= 'b0;
		  data <= 'b0;
        $readmemh("/home/alejandro/github-classroom/digital-electronics-UNAL/lab07-lcd-en-modo-paralelo-2025-ii-ed-g5-e1/src/data.txt", static_data_mem);
    end else begin
        case (next_state)
            IDLE: begin
                command_counter <= 'b0;
                data_counter <= 'b0;
                rs <= 1'b0;
                data  <= 'b0;
            end
            CONFIG_CMD1: begin
			    rs <= 1'b0; 	
                command_counter <= command_counter + 1;
				data <= config_mem[command_counter];
            end
            WR_STATIC_TEXT_1L: begin
                data_counter <= data_counter + 1;
                rs <= 1'b1; 
				data <= static_data_mem[data_counter];
            end
            CONFIG_CMD2: begin
                data_counter <= 'b0;
				rs <= 1'b0; 
				data <= START_2LINE;
            end
			WR_STATIC_TEXT_2L: begin
                data_counter <= data_counter + 1;
                rs <= 1'b1; 
				data <= static_data_mem[NUM_DATA_PERLINE + data_counter];
            end
        endcase
    end
end

assign enable = clk_16ms;

endmodule
